module gw_gao(
    \uart_rx_bytes[23] ,
    \uart_rx_bytes[22] ,
    \uart_rx_bytes[21] ,
    \uart_rx_bytes[20] ,
    \uart_rx_bytes[19] ,
    \uart_rx_bytes[18] ,
    \uart_rx_bytes[17] ,
    \uart_rx_bytes[16] ,
    \uart_rx_bytes[15] ,
    \uart_rx_bytes[14] ,
    \uart_rx_bytes[13] ,
    \uart_rx_bytes[12] ,
    \uart_rx_bytes[11] ,
    \uart_rx_bytes[10] ,
    \uart_rx_bytes[9] ,
    \uart_rx_bytes[8] ,
    \uart_rx_bytes[7] ,
    \uart_rx_bytes[6] ,
    \uart_rx_bytes[5] ,
    \uart_rx_bytes[4] ,
    \uart_rx_bytes[3] ,
    \uart_rx_bytes[2] ,
    \uart_rx_bytes[1] ,
    \uart_rx_bytes[0] ,
    clk,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input \uart_rx_bytes[23] ;
input \uart_rx_bytes[22] ;
input \uart_rx_bytes[21] ;
input \uart_rx_bytes[20] ;
input \uart_rx_bytes[19] ;
input \uart_rx_bytes[18] ;
input \uart_rx_bytes[17] ;
input \uart_rx_bytes[16] ;
input \uart_rx_bytes[15] ;
input \uart_rx_bytes[14] ;
input \uart_rx_bytes[13] ;
input \uart_rx_bytes[12] ;
input \uart_rx_bytes[11] ;
input \uart_rx_bytes[10] ;
input \uart_rx_bytes[9] ;
input \uart_rx_bytes[8] ;
input \uart_rx_bytes[7] ;
input \uart_rx_bytes[6] ;
input \uart_rx_bytes[5] ;
input \uart_rx_bytes[4] ;
input \uart_rx_bytes[3] ;
input \uart_rx_bytes[2] ;
input \uart_rx_bytes[1] ;
input \uart_rx_bytes[0] ;
input clk;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire \uart_rx_bytes[23] ;
wire \uart_rx_bytes[22] ;
wire \uart_rx_bytes[21] ;
wire \uart_rx_bytes[20] ;
wire \uart_rx_bytes[19] ;
wire \uart_rx_bytes[18] ;
wire \uart_rx_bytes[17] ;
wire \uart_rx_bytes[16] ;
wire \uart_rx_bytes[15] ;
wire \uart_rx_bytes[14] ;
wire \uart_rx_bytes[13] ;
wire \uart_rx_bytes[12] ;
wire \uart_rx_bytes[11] ;
wire \uart_rx_bytes[10] ;
wire \uart_rx_bytes[9] ;
wire \uart_rx_bytes[8] ;
wire \uart_rx_bytes[7] ;
wire \uart_rx_bytes[6] ;
wire \uart_rx_bytes[5] ;
wire \uart_rx_bytes[4] ;
wire \uart_rx_bytes[3] ;
wire \uart_rx_bytes[2] ;
wire \uart_rx_bytes[1] ;
wire \uart_rx_bytes[0] ;
wire clk;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(1'b0)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top u_ao_top(
    .control(control0[9:0]),
    .data_i({\uart_rx_bytes[23] ,\uart_rx_bytes[22] ,\uart_rx_bytes[21] ,\uart_rx_bytes[20] ,\uart_rx_bytes[19] ,\uart_rx_bytes[18] ,\uart_rx_bytes[17] ,\uart_rx_bytes[16] ,\uart_rx_bytes[15] ,\uart_rx_bytes[14] ,\uart_rx_bytes[13] ,\uart_rx_bytes[12] ,\uart_rx_bytes[11] ,\uart_rx_bytes[10] ,\uart_rx_bytes[9] ,\uart_rx_bytes[8] ,\uart_rx_bytes[7] ,\uart_rx_bytes[6] ,\uart_rx_bytes[5] ,\uart_rx_bytes[4] ,\uart_rx_bytes[3] ,\uart_rx_bytes[2] ,\uart_rx_bytes[1] ,\uart_rx_bytes[0] }),
    .clk_i(clk)
);

endmodule
